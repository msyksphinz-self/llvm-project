assign A = 0;
assign Hoge = A;
