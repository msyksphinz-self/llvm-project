assign A = 3;
assign B = 4;

assign Hoge1 = A + B;
assign Hoge2 = A * B;
