assign A = 0;
assign Hoge = 2;
