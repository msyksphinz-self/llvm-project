assign A = 3;
assign Hoge = A;
assign B = 4;
assign Hoge = B;
